hihhbhjhb
